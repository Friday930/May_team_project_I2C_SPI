`timescale 1ns / 1ps

module SPI_Master (
    input            clk,
    input            reset,
    input            cpol,     //새로이 추가된
    input            cpha,     // 상태에 따른 clk변화
    input            start,
    input   ss, // 수정 부분***
    output     [7:0] rx_data,
    input      [7:0] tx_data,
    output reg       done,
    output reg       ready,
    output           SCLK,
    output           MOSI,
    input            MISO,
    output SS // 수정 부분***
);
    parameter IDLE = 0, CP_DELAY = 1, CP0 = 2, CP1 = 3;

    wire r_sclk;
    reg [1:0] state, state_next;
    reg [7:0] temp_tx_data_reg, temp_tx_data_next;
    reg [7:0] temp_rx_data_reg, temp_rx_data_next;
    reg [5:0] sclk_counter_reg, sclk_counter_next;
    reg [2:0] bit_counter_reg, bit_counter_next;

    assign SS = ss;
    assign MOSI = temp_tx_data_reg[7];
    assign rx_data = temp_rx_data_reg;

    assign r_sclk = (state_next == CP1 && ~cpha) || (state_next == CP0 && cpha);
    // r_sclk가 high 출력이 되는 조건 -> CPOL이 0일 때
    assign SCLK = cpol ? ~r_sclk : r_sclk; // CPOL이 1이면 반전 0이면 유지

    always @(posedge clk, posedge reset) begin
        if (reset) begin
            state <= IDLE;
            temp_tx_data_reg <= 0;
            temp_rx_data_reg <= 8'd0;
            sclk_counter_reg <= 0;
            bit_counter_reg <= 0;
        end else begin
            state <= state_next;
            temp_tx_data_reg <= temp_tx_data_next;
            temp_rx_data_reg <= temp_rx_data_next;
            sclk_counter_reg <= sclk_counter_next;
            bit_counter_reg <= bit_counter_next;
        end
    end

    always @(*) begin
        state_next        = state;
        done              = 0;
        ready             = 0;
        
        temp_rx_data_next = temp_rx_data_reg;
        temp_tx_data_next = temp_tx_data_reg;
        sclk_counter_next = sclk_counter_reg;
        bit_counter_next  = bit_counter_reg;
        case (state)
            IDLE: begin
                temp_tx_data_next = 0;
                done = 0;
                ready = 1;
                if (start) begin
                    state_next = cpha ? CP_DELAY : CP0; //CPHA에따라서 0과 1일때의 차이는 CP0가 나타나기 전 DELAY 발생 여부
                    temp_tx_data_next = tx_data;
                    ready = 0;
                    sclk_counter_next = 0;
                    bit_counter_next = 0;
                end
            end
            CP_DELAY: begin
                if (sclk_counter_reg == 49) begin
                    sclk_counter_next = 0;
                    state_next = CP0;
                end else begin
                    sclk_counter_next = sclk_counter_reg + 1;
                end
            end
            CP0: begin
                //r_sclk = 0;
                if (sclk_counter_reg == 49) begin
                    temp_rx_data_next = {temp_rx_data_reg[6:0], MISO};
                    sclk_counter_next = 0;
                    state_next = CP1;
                end else begin
                    sclk_counter_next = sclk_counter_reg + 1;
                end
            end
            CP1: begin
                //r_sclk = 1'b1;
                if (sclk_counter_reg == 49) begin
                    if (bit_counter_reg == 7) begin
                        state_next = IDLE;
                        done = 1'b1;
                    end else begin
                        temp_tx_data_next = {temp_tx_data_reg[6:0], 1'b0};
                        sclk_counter_next = 6'd0;
                        bit_counter_next = bit_counter_reg + 1;
                        state_next = CP0;
                    end
                end else begin
                    sclk_counter_next = sclk_counter_reg + 1;
                end
            end
        endcase
    end
endmodule
